module cla_32_gen(input [31:0]a,input [31:0]b,input carry_in,output [31:0]c);


wire  [31:0]p,g;


assign p[0]=a[0]^b[0];
assign g[0]=a[0]&b[0];
assign p[1]=a[1]^b[1];
assign g[1]=a[1]&b[1];
assign p[2]=a[2]^b[2];
assign g[2]=a[2]&b[2];
assign p[3]=a[3]^b[3];
assign g[3]=a[3]&b[3];

assign p[4]=a[4]^b[4];
assign g[4]=a[4]&b[4];
assign p[5]=a[5]^b[5];
assign g[5]=a[5]&b[5];
assign p[6]=a[6]^b[6];
assign g[6]=a[6]&b[6];
assign p[7]=a[7]^b[7];
assign g[7]=a[7]&b[7];
assign p[8]=a[8]^b[8];
assign g[8]=a[8]&b[8];
assign p[9]=a[9]^b[9];
assign g[9]=a[9]&b[9];
assign p[10]=a[10]^b[10];
assign g[10]=a[10]&b[10];
assign p[11]=a[11]^b[11];
assign g[11]=a[11]&b[11];
assign p[12]=a[12]^b[12];
assign g[12]=a[12]&b[12];
assign p[13]=a[13]^b[13];
assign g[13]=a[13]&b[13];
assign p[14]=a[14]^b[14];
assign g[14]=a[14]&b[14];
assign p[15]=a[15]^b[15];
assign g[15]=a[15]&b[15];
assign p[16]=a[16]^b[16];
assign g[16]=a[16]&b[16];
assign p[17]=a[17]^b[17];
assign g[17]=a[17]&b[17];
assign p[18]=a[18]^b[18];
assign g[18]=a[18]&b[18];
assign p[19]=a[19]^b[19];
assign g[19]=a[19]&b[19];
assign p[20]=a[20]^b[20];
assign g[20]=a[20]&b[20];
assign p[21]=a[21]^b[21];
assign g[21]=a[21]&b[21];
assign p[22]=a[22]^b[22];
assign g[22]=a[22]&b[22];
assign p[23]=a[23]^b[23];
assign g[23]=a[23]&b[23];
assign p[24]=a[24]^b[24];
assign g[24]=a[24]&b[24];
assign p[25]=a[25]^b[25];
assign g[25]=a[25]&b[25];
assign p[26]=a[26]^b[26];
assign g[26]=a[26]&b[26];
assign p[27]=a[27]^b[27];
assign g[27]=a[27]&b[27];
assign p[28]=a[28]^b[28];
assign g[28]=a[28]&b[28];
assign p[29]=a[29]^b[29];
assign g[29]=a[29]&b[29];
assign p[30]=a[30]^b[30];
assign g[30]=a[30]&b[30];
assign p[31]=a[31]^b[31];
assign g[31]=a[31]&b[31];



assign c[0]=(p[0] & carry_in) | g[0];
assign c[1]=(p[1] & p[0] & carry_in)|(p[1] & g[0]) | g[1];
assign c[2]=(p[2] & p[1] & p[0] & carry_in)|(p[2] & p[1] & g[0]) | (p[2] & g[1]) | g[2];
assign c[3]=(p[3] & p[2] & p[1] & p[0] & carry_in)|(p[3] & p[2] & p[1] & g[0])|(p[3] & p[2] & g[1]) | (p[3] & g[2]) | g[3];

assign c[4]=(p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[4]&p[3]&p[2]&p[1]&g[0])|(p[4]&p[3]&p[2]&g[1])|(p[4]&p[3]&g[2])|(p[4]&g[3])|g[4];
assign c[5]=(p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[5]&p[4]&p[3]&p[2]&g[1])|(p[5]&p[4]&p[3]&g[2])|(p[5]&p[4]&g[3])|(p[5]&g[4])|g[5];
assign c[6]=(p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[6]&p[5]&p[4]&p[3]&g[2])|(p[6]&p[5]&p[4]&g[3])|(p[6]&p[5]&g[4])|(p[6]&g[5])|(g[6]);
assign c[7]=(p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[7]&p[6]&p[5]&p[4]&g[3])|(p[7]&p[6]&p[5]&g[4])|(p[7]&p[6]&g[5])|(p[7]&g[6])|(g[7]);
assign c[8]=(p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[8]&p[7]&p[6]&p[5]&g[4])|(p[8]&p[7]&p[6]&g[5])|(p[8]&p[7]&g[6])|(p[8]&g[7])|(g[8]);
assign c[9]=(p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[9]&p[8]&p[7]&p[6]&g[5])|(p[9]&p[8]&p[7]&g[6])|(p[9]&p[8]&g[7])|(p[9]&g[8])|(g[9]);
assign c[10]=(p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[10]&p[9]&p[8]&p[7]&g[6])|(p[10]&p[9]&p[8]&g[7])|(p[10]&p[9]&g[8])|(p[10]&g[9])|(g[10]);

assign c[11]=(p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[11]&p[10]&p[9]&p[8]&g[7])|(p[11]&p[10]&p[9]&g[8])|(p[11]&p[10]&g[9])|(p[11]&g[10])|(g[11]);
assign c[12]=(p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[12]&p[11]&p[10]&p[9]&g[8])|(p[12]&p[11]&p[10]&g[9])|(p[12]&p[11]&g[10])|(p[12]&g[11])|(g[12]);
assign c[13]=(p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[13]&p[12]&p[11]&p[10]&g[9])|(p[13]&p[12]&p[11]&g[10])|(p[13]&p[12]&g[11])|(p[13]&g[12])|(g[13]);
assign c[14]=(p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[14]&p[13]&p[12]&p[11]&p[10]&g[9])|(p[14]&p[13]&p[12]&p[11]&g[10])|(p[14]&p[13]&p[12]&g[11])|(p[14]&p[13]&g[12])|(p[14]&g[13])|(g[14]);
assign c[15]=(p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9])|(p[15]&p[14]&p[13]&p[12]&p[11]&g[10])|(p[15]&p[14]&p[13]&p[12]&g[11])|(p[15]&p[14]&p[13]&g[12])|(p[15]&p[14]&g[13])|(p[15]&g[14])|(g[15]);
assign c[16]=(p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9])|(p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&g[10])|(p[16]&p[15]&p[14]&p[13]&p[12]&g[11])|(p[16]&p[15]&p[14]&p[13]&g[12])|(p[16]&p[15]&p[14]&g[13])|(p[16]&p[15]&g[14])|(p[16]&g[15])|(g[16]);
assign c[17]=(p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9])|(p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&g[10])|(p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&g[11])|(p[17]&p[16]&p[15]&p[14]&p[13]&g[12])|(p[17]&p[16]&p[15]&p[14]&g[13])|(p[17]&p[16]&p[15]&g[14])|(p[17]&p[16]&g[15])|(p[17]&g[16])|(g[17]);
assign c[18]=(p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9])|(p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&g[10])|(p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&g[11])|(p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&g[12])|(p[18]&p[17]&p[16]&p[15]&p[14]&g[13])|(p[18]&p[17]&p[16]&p[15]&g[14])|(p[18]&p[17]&p[16]&g[15])|(p[18]&p[17]&g[16])|(p[18]&g[17])|(g[18]);
assign c[19]=(p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9])|(p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&g[10])|(p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&g[11])|(p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&g[12])|(p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&g[13])|(p[19]&p[18]&p[17]&p[16]&p[15]&g[14])|(p[19]&p[18]&p[17]&p[16]&g[15])|(p[19]&p[18]&p[17]&g[16])|(p[19]&p[18]&g[17])|(p[19]&g[18])|(g[19]);
assign c[20]=(p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9])|(p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&g[10])|(p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&g[11])|(p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&g[12])|(p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&g[13])|(p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&g[14])|(p[20]&p[19]&p[18]&p[17]&p[16]&g[15])|(p[20]&p[19]&p[18]&p[17]&g[16])|(p[20]&p[19]&p[18]&g[17])|(p[20]&p[19]&g[18])|(p[20]&g[19])|g[20];
assign c[21]=(p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9])|(p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&g[10])|(p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&g[11])|(p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&g[12])|(p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&g[13])|(p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&g[14])|(p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&g[15])|(p[21]&p[20]&p[19]&p[18]&p[17]&g[16])|(p[21]&p[20]&p[19]&p[18]&g[17])|(p[21]&p[20]&p[19]&g[18])|(p[21]&p[20]&g[19])|(p[21]&g[20])|(g[21]);
assign c[22]=(p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9])|(p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&g[10])|(p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&g[11])|(p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&g[12])|(p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&g[13])|(p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&g[14])|(p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&g[15])|(p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&g[16])|(p[22]&p[21]&p[20]&p[19]&p[18]&g[17])|(p[22]&p[21]&p[20]&p[19]&g[18])|(p[22]&p[21]&p[20]&g[19])|(p[22]&p[21]&g[20])|(p[22]&g[21])|(g[22]);
assign c[23]=(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9])|(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&g[10])|(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&g[11])|(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&g[12])|(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&g[13])|(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&g[14])|(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&g[15])|(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&g[16])|(p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&g[17])|(p[23]&p[22]&p[21]&p[20]&p[19]&g[18])|(p[23]&p[22]&p[21]&p[20]&g[19])|(p[23]&p[22]&p[21]&g[20])|(p[23]&p[22]&g[21])|(p[23]&g[22])|(g[23]);
assign c[24]=(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9])|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&g[10])|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&g[11])|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&g[12])|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&g[13])|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&g[14])|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&g[15])|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&g[16])|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&g[17])|(p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&g[18])|(p[24]&p[23]&p[22]&p[21]&p[20]&g[19])|(p[24]&p[23]&p[22]&p[21]&g[20])|(p[24]&p[23]&p[22]&g[21])|(p[24]&p[23]&g[22])|(p[24]&g[23])|(g[24]);
assign c[25]=(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&g[10])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&g[11])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&g[12])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&g[13])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&g[14])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&g[15])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&g[16])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&g[17])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&g[18])|(p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&g[19])|(p[25]&p[24]&p[23]&p[22]&p[21]&g[20])|(p[25]&p[24]&p[23]&p[22]&g[21])|(p[25]&p[24]&p[23]&g[22])|(p[25]&p[24]&g[23])|(p[25]&p[24]&g[23])|(p[25]&g[24])|(g[25]);
assign c[26]=(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&g[10])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&g[11])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&g[12])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&g[13])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&g[14])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&g[15])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&g[16])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&g[17])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&g[18])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&g[19])|(p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&g[20])|(p[26]&p[25]&p[24]&p[23]&p[22]&g[21])|(p[26]&p[25]&p[24]&p[23]&g[22])|(p[26]&p[25]&p[24]&g[23])|(p[26]&p[25]&p[24]&g[23])|(p[26]&p[25]&g[24])|(p[26]&g[25])|(g[26]);
assign c[27]=(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&g[10])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&g[11])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&g[12])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&g[13])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&g[14])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&g[15])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&g[16])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&g[17])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&g[18])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&g[19])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&g[20])|(p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&g[21])|(p[27]&p[26]&p[25]&p[24]&p[23]&g[22])|(p[27]&p[26]&p[25]&p[24]&g[23])|(p[27]&p[26]&p[25]&p[24]&g[23])|(p[27]&p[26]&p[25]&g[24])|(p[27]&p[26]&g[25])|(p[27]&g[26])|(g[27]);
assign c[28]=(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&g[10])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&g[11])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&g[12])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&g[13])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&g[14])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&g[15])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&g[16])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&g[17])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&g[18])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&g[19])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&g[20])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&g[21])|(p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&g[22])|(p[28]&p[27]&p[26]&p[25]&p[24]&g[23])|(p[28]&p[27]&p[26]&p[25]&p[24]&g[23])|(p[28]&p[27]&p[26]&p[25]&g[24])|(p[28]&p[27]&p[26]&g[25])|(p[28]&p[27]&g[26])|(p[28]&g[27])|(g[28]);
assign c[29]=(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&g[10])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&g[11])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&g[12])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&g[13])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&g[14])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&g[15])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&g[16])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&g[17])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&g[18])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&g[19])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&g[20])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&g[21])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&g[22])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&g[23])|(p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&g[23])|(p[29]&p[28]&p[27]&p[26]&p[25]&g[24])|(p[29]&p[28]&p[27]&p[26]&g[25])|(p[29]&p[28]&p[27]&g[26])|(p[29]&p[28]&g[27])|(p[29]&g[28])|(g[29]);
assign c[30]=(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&g[10])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&g[11])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&g[12])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&g[13])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&g[14])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&g[15])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&g[16])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&g[17])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&g[18])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&g[19])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&g[20])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&g[21])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&g[22])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&g[23])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&g[23])|(p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&g[24])|(p[30]&p[29]&p[28]&p[27]&p[26]&g[25])|(p[30]&p[29]&p[28]&p[27]&g[26])|(p[30]&p[29]&p[28]&g[27])|(p[30]&p[29]&g[28])|(p[30]&g[29])|(g[30]);
assign c[31]=(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&p[0]&carry_in)|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&p[1]&g[0])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&p[2]&g[1])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&p[3]&g[2])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&p[4]&g[3])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&p[5]&g[4])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&p[6]&g[5])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&p[7]&g[6])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&p[8]&g[7])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&p[9]&g[8])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&p[10]&g[9])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&p[11]&g[10])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&p[12]&g[11])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&p[13]&g[12])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&p[14]&g[13])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&p[15]&g[14])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&p[16]&g[15])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&p[17]&g[16])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&p[18]&g[17])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&p[19]&g[18])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&p[20]&g[19])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&p[21]&g[20])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&p[22]&g[21])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&p[23]&g[22])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&g[23])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&p[24]&g[23])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&p[25]&g[24])|(p[31]&p[30]&p[29]&p[28]&p[27]&p[26]&g[25])|(p[31]&p[30]&p[29]&p[28]&p[27]&g[26])|(p[31]&p[30]&p[29]&p[28]&g[27])|(p[31]&p[30]&p[29]&g[28])|(p[31]&p[30]&g[29])|(p[31]&g[30])|(g[31]);

 

endmodule